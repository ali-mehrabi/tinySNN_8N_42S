module neucleus
(parameter p_width = 8);
(
input   [p_width-1:0]  i_a,
input   [p_width-1:0]  i_b,
input   [p_width-1:0]  i_c,
input   [p_width-1:0]  i_d,
output                 o_s
); 




endmodule